`timescale 1ns / 1ps
/////////////////////////////////////
module hw1(
    );


endmodule
